// uart.vh

`define IDLE_BIT  1'b1
`define START_BIT 1'b0
`define STOP_BIT  1'b1
